/***********************************************************************
 * A SystemVerilog testbench for an instruction register.
 * The course labs will convert this to an object-oriented testbench
 * with constrained random test generation, functional coverage, and
 * a scoreboard for self-verification.
 **********************************************************************/

module instr_register_test
  import instr_register_pkg::*;  // user-defined types are defined in instr_register_pkg.sv
(
    input  logic         clk,
    output logic         load_en,
    output logic         reset_n,
    output operand_t     operand_a,
    output operand_t     operand_b,
    output opcode_t      opcode,
    output address_t     write_pointer,
    output address_t     read_pointer,
    input  instruction_t instruction_word
);

  timeunit 1ns / 1ns;
  parameter read_number = 20, write_number = 20;
  int number_of_errors_per_test = 0;
  int seed = 555;

  initial begin
    $display("\n\n***********************************************************");
    $display("***  THIS IS NOT A SELF-CHECKING TESTBENCH (YET).  YOU  ***");
    $display("***  NEED TO VISUALLY VERIFY THAT THE OUTPUT VALUES     ***");
    $display("***  MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display("***********************************************************");

    $display("\nReseting the instruction register...");
    write_pointer = 5'h00;  // initialize write pointer
    read_pointer  = 5'h1F;  // initialize read pointer
    load_en       = 1'b0;  // initialize load control line
    reset_n <= 1'b0;  // assert reset_n (active low)
    repeat (2) @(posedge clk);  // hold in reset for 2 clock cycles
    reset_n = 1'b1;  // deassert reset_n (active low)

    $display("\nWriting values to register stack...");
    @(posedge clk) load_en = 1'b1;  // enable writing to register
    // A.M. 9:19 - 11/3/2024 
    //repeat (3) begin
    repeat (write_number) begin
      @(posedge clk) randomize_transaction;
      @(negedge clk) print_transaction;
    end
    @(posedge clk) load_en = 1'b0;  // turn-off writing to register

    // read back and display same three register locations
    $display("\nReading back the same register locations written...");
    // A.M. 9:19 - 11/3/2024 
    // for (int i=0; i<=2; i++) begin
    for (int i = 0; i <= read_number; i++) begin
      // later labs will replace this loop with iterating through a
      // scoreboard to determine which addresses were written and
      // the expected values to be read back
      @(posedge clk) read_pointer = i;
      @(negedge clk) print_results;
      check_result;
    end

    @(posedge clk);
    $display("\nNumber of errors during TEST: %0d", number_of_errors_per_test);
    $display("\n***********************************************************");
    $display("***  THIS IS NOT A SELF-CHECKING TESTBENCH (YET).  YOU  ***");
    $display("***  NEED TO VISUALLY VERIFY THAT THE OUTPUT VALUES     ***");
    $display("***  MATCH THE INPUT VALUES FOR EACH REGISTER LOCATION  ***");
    $display("***********************************************************\n");
    $finish;
  end

  function void randomize_transaction;
    // A later lab will replace this function with SystemVerilog
    // constrained random values
    //
    // The stactic temp variable is required in order to write to fixed
    // addresses of 0, 1 and 2.  This will be replaceed with randomizeed
    // write_pointer values in a later lab
    //
    static int temp = 0;
    operand_a     <= $random(seed) % 16;  // between -15 and 15
    operand_b     <= $unsigned($random) % 16;  // between 0 and 15
    opcode        <= opcode_t'($unsigned($random) % 8);  // between 0 and 7, cast to opcode_t type
    write_pointer <= temp++;
  endfunction : randomize_transaction

  function void print_transaction;
    $display("Writing to register location %0d: ", write_pointer);
    $display("  opcode = %0d (%s)", opcode, opcode.name);
    $display("  operand_a = %0d", operand_a);
    $display("  operand_b = %0d\n", operand_b);
  endfunction : print_transaction

  function void print_results;
    $display("Read from register location %0d: ", read_pointer);
    $display("  opcode = %0d (%s)", instruction_word.opc, instruction_word.opc.name);
    $display("  operand_a = %0d", instruction_word.op_a);
    $display("  operand_b = %0d", instruction_word.op_b);
    $display("  result = %0d\n", instruction_word.result);
  endfunction : print_results

  function void check_result;
    operand_result_t exp_result;

    if (instruction_word.opc == ZERO) begin
      exp_result = 'b0;
    end else if (instruction_word.opc == PASSA) begin
      exp_result = instruction_word.op_a;
    end else if (instruction_word.opc == PASSB) begin
      exp_result = instruction_word.op_b;
    end else if (instruction_word.opc == ADD) begin
      exp_result = instruction_word.op_a + instruction_word.op_b;
    end else if (instruction_word.opc == SUB) begin
      exp_result = instruction_word.op_a - instruction_word.op_b;
    end else if (instruction_word.opc == MULT) begin
      exp_result = instruction_word.op_a * instruction_word.op_b;
    end else if (instruction_word.opc == DIV) begin
      if (instruction_word.op_b == 0) begin
        number_of_errors_per_test++;
        return;
      end else begin
        exp_result = instruction_word.op_a / instruction_word.op_b;
      end
    end else if (instruction_word.opc == MOD) begin
      exp_result = instruction_word.op_a % instruction_word.op_b;
    end

    if (exp_result != instruction_word.result) begin
      number_of_errors_per_test++;
    end
  endfunction : check_result
endmodule : instr_register_test
